package lab;
module lab ();
    rule main;
        $display("Hello, world!");
        $finish();
    endrule
endmodule
endpackage